



`timescale 1ns / 1ps 

// RANDOM GOLDEN SELF CHECKING TEST BENCH,  
// This test bench generates random single instructions (not a sequence)
// resets the processor, initializes instruction memory and data memory
// randomly and then runs the processor to execute the instructon checking if
// the processor is executing the instruction correctly or not. 
// // // // // 



module riscv32isinglecycle_singleInstruction_rand_tb(); 

reg clk; 
reg rst;












endmodule
